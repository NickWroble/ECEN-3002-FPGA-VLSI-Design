
module ISSP_KEY (
	source,
	probe);	

	output	[2:0]	source;
	input	[2:0]	probe;
endmodule
